module bch (s, d);
input [3:0] s;
output reg [6:0] d;

always @(s)
case({s})
	4'b0000 : d<= 7'b1000000;
	4'b0001 : d<= 7'b1111001;
	4'b0010 : d<= 7'b0100100;
	4'b0011 : d<= 7'b0110000;
	4'b0100 : d<= 7'b0011001;
	4'b0101 : d<= 7'b0010010;
	4'b0110 : d<= 7'b0000010;
	4'b0111 : d<= 7'b1111000;
	4'b1000 : d<= 7'b0000000;
	4'b1001 : d<= 7'b0011000;
	4'b1010 : d<= 7'b0001000;
	4'b1011 : d<= 7'b0000011;
	4'b1100 : d<= 7'b1000110;
	4'b1101 : d<= 7'b0100001;
	4'b1110 : d<= 7'b0000110;
	4'b1111 : d<= 7'b0001110;	
endcase	
endmodule 